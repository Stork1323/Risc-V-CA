module Stage_Ex( // stage execute 
	input logic [31:0] R1_i, R2_i,
	output logic [31:0] A_o, B_o
	);
	
	
	
endmodule
