module Stage_Mem( // stage memory access
	);
	
endmodule
