`ifndef DEFINE_sv
`define DEFINE_sv

`define OP_Rtype 		 0110011
`define OP_Itype 		 0010011
`define OP_Itype_load 0000011
`define OP_Stype 		 0100011
`define OP_Btype 		 1100011
`define OP_JAL 		 1101111
`define OP_LUI 		 0110111
`define OP_AUIPC 		 0010111
`define OP_JALR 		 1100111



`endif
