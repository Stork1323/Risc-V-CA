module Stage_Wb( // stage write back to register
	);
	
endmodule

